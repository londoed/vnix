module file
