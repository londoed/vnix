module main

import asm
import dev
import fs
import lock
import mem
import proc
import sys
