module dev

import asm
import fs
import lock
import mem
import proc
import sys
