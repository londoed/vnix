module syscall

import types
import defs
import param
import memlay
import mmu
import proc
import x86
import syscall
