module asm

// NEED INLINE ASSEMBLER!
