module types

pub type pde_t byte
