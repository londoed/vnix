module vnix

pub type pde_t byte
