module sys

pub struct RTCDate {
pub mut:
	second u32
	minute u32
	hour u32
	day u32
	month u32
	year u32
}
